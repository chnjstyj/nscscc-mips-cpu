module mem(
    input [31:0] ALU_result,
    input [31:0] din,
    input MemWrite,
    input MemRead,
    input MemtoReg,
    output [31:0] dout
);




endmodule 