module top(
    input clk,
    input rst
);

wire ce;
wire [31:0] inst_address;
wire [31:0] cur_inst;
wire [31:0] next_instaddress;
wire [5:0] opcode;
wire [4:0] rreg_a;
wire [4:0] rreg_b;
wire [4:0] wreg;
wire [31:0] imme_num;
wire [5:0] func;
wire [3:0] alu_control_sig;
wire ALU_zerotag;
wire [4:0] shamt;
wire bgtz_sig;

//id�׶ο����ź�
wire RegDst;
wire Branch;
wire MemRead;
wire MemtoReg;
wire [3:0] ALUOp;
wire MemWrite;
wire ALUSrc;
wire RegWrite;
wire Jump;                    //�͵�ƽ��Ч
wire unsigned_num;           //��ʱ����
wire equal_branch;
wire store_pc;
wire lui_sig;
wire greater_than;
wire zero_sig;

//ex�׶ο����ź�
wire jmp_reg;                //jr �ź���

//��ַ������
wire [31:0] jc_instaddress;

//�Ĵ����Ѷ�������
wire [31:0] rdata_a;
wire [31:0] rdata_b;

//alu����
wire [31:0] alu_rdata_a;
wire [31:0] alu_rdata_b;

//alu������
wire [31:0] alu_result;

//������Ƭѡ�ź�
wire [1:0] mem_sel;

//�������������� //�Ĵ���д���ַ �Ĵ���д���ź�
wire [31:0] mem_wdata;
/*wire [4:0] wb_wreg;
wire wb_RegWrite;*/

//��·�������
wire control_rdata_a;
wire control_rdata_b;

//��ˮ������ģ������
wire stall_if_id;
wire stall_id_ex;
wire stall_ex_memwb;

//��ˮ�����ģ��������
//if_id
wire [31:0] id_inst;
wire [31:0] id_next_instaddress;
wire [31:0] id_cur_instaddress;
if_id if_id(
    .clk(clk),
    .rst(rst),
    .if_inst(cur_inst),
    .if_next_instaddress(next_instaddress),
    .if_cur_instaddress(inst_address),
    .stall_if_id(stall_if_id),
    .id_inst(id_inst),
    .id_next_instaddress(id_next_instaddress),
    .id_cur_instaddress(id_cur_instaddress)
);

//id_ex
wire ex_Branch;
wire ex_MemRead;
wire ex_MemtoReg;
wire [3:0] ex_ALUOp;
wire ex_MemWrite;
wire ex_ALUSrc;
wire ex_RegWrite;
wire ex_equal_branch;
wire ex_lui_sig;
wire [31:0] ex_next_instaddress;
wire [31:0] ex_rdata_a;
wire [31:0] ex_rdata_b;
wire [31:0] ex_imme_num;
wire [5:0] ex_func;
wire [4:0] ex_shamt;
wire [5:0] ex_opcode;
wire [31:0] ex_cur_instaddress;
wire [4:0] ex_wreg;
wire [4:0] ex_Rs;
wire [4:0] ex_Rt;
wire ex_greater_than;
 
id_ex id_ex(
    .clk(clk),
    .rst(rst),
    .stall_id_ex(stall_id_ex),
    //.id_Branch(Branch),
    .id_MemRead(MemRead),
    .id_MemtoReg(MemtoReg),
    .id_ALUOp(ALUOp),
    .id_MemWrite(MemWrite),
    .id_ALUSrc(ALUSrc),
    .id_RegWrite(RegWrite),
    .id_equal_branch(equal_branch),
    .id_store_pc(store_pc),
    .id_lui_sig(lui_sig),
    .id_next_instaddress(id_next_instaddress),
    .id_rdata_a(rdata_a),
    .id_rdata_b(rdata_b),
    .id_imme_num(imme_num),
    .id_func(func),
    .id_shamt(shamt),
    .id_opcode(opcode),
    .id_cur_instaddress(id_cur_instaddress),
    .id_wreg(wreg),
    .id_Rs(rreg_a),
    .id_Rt(rreg_b),
    .id_greater_than(greater_than),
   // .ex_Branch(ex_Branch),
    .ex_MemRead(ex_MemRead),
    .ex_MemtoReg(ex_MemtoReg),
    .ex_ALUOp(ex_ALUOp),
    .ex_MemWrite(ex_MemWrite),
    .ex_ALUSrc(ex_ALUSrc),
    .ex_RegWrite(ex_RegWrite),
    .ex_equal_branch(ex_equal_branch),
    .ex_store_pc(ex_store_pc),
    .ex_lui_sig(ex_lui_sig),
    .ex_next_instaddress(ex_next_instaddress),
    .ex_rdata_a(ex_rdata_a),
    .ex_rdata_b(ex_rdata_b),
    .ex_imme_num(ex_imme_num),
    .ex_func(ex_func),
    .ex_shamt(ex_shamt),
    .ex_opcode(ex_opcode),
    .ex_cur_instaddress(ex_cur_instaddress),
    .ex_wreg(ex_wreg),
    .ex_Rs(ex_Rs),
    .ex_Rt(ex_Rt),
    .ex_greater_than(ex_greater_than)
);

//ex_mem
wire mem_lui_sig;
wire mem_MemRead;
wire mem_MemWrite;
wire mem_MemtoReg;
wire mem_RegWrite;
wire [31:0] mem_alu_result;
wire [31:0] mem_rdata_b;
wire [5:0] mem_opcode;
wire [31:0] mem_imme_num;
wire [4:0] mem_wreg;
ex_mem ex_mem(
    .clk(clk),
    .rst(rst),
    .ex_lui_sig(ex_lui_sig),
    .ex_MemRead(ex_MemRead),
    .ex_MemWrite(ex_MemWrite),
    .ex_MemtoReg(ex_MemtoReg),
    .ex_RegWrite(ex_RegWrite),
    .ex_alu_result(alu_result),
    .ex_rdata_b(ex_rdata_b),
    .ex_opcode(ex_opcode),
    .ex_imme_num(ex_imme_num),
    .ex_wreg(ex_wreg),
    .mem_lui_sig(mem_lui_sig),
    .mem_MemRead(mem_MemRead),
    .mem_MemWrite(mem_MemWrite),
    .mem_MemtoReg(mem_MemtoReg),
    .mem_RegWrite(mem_RegWrite),
    .mem_alu_result(mem_alu_result),
    .mem_rdata_b(mem_rdata_b),
    .mem_opcode(mem_opcode),
    .mem_imme_num(mem_imme_num),
    .mem_wreg(mem_wreg)
);

//��ˮ������ģ��
stall stall(
    .Jump(Jump),
    .jmp_reg(jmp_reg),
    .id_Branch(Branch),
    .zero_sig(zero_sig),
    .bgtz_sig(bgtz_sig),
    .stall_if_id(stall_if_id),
    .stall_id_ex(stall_id_ex),
    .stall_ex_memwb(stall_ex_memwb)
);

pc pc(
    .clk(clk),
    .rst(rst),
    .Branch(Branch),
    .zero_sig(zero_sig),
    .Jump(Jump),
    .imme(imme_num),
    .jmp_reg(jmp_reg),
    .Rrs(ex_rdata_a),                
    .jc_instaddress(jc_instaddress),
    .id_cur_inst(id_inst),
    .id_next_instaddress(id_next_instaddress),
    .inst_address(inst_address),
    .next_instaddress(next_instaddress),
    .bgtz_sig(bgtz_sig),
    .ce(ce)
);

inst_reg inst_reg(
    .clk(clk),
    .inst_address(inst_address),
    .ce(ce),
    .inst(cur_inst)
);

id id(
    .inst(id_inst),
    .RegDst(RegDst),
    .opcode(opcode),
    .rreg_a(rreg_a),
    .rreg_b(rreg_b),
    .wreg(wreg),
    .imme_num(imme_num),
    .func(func),
    .shamt(shamt),
    .jmp_reg
);

branch branch(
    .next_instaddress(id_next_instaddress),          //����id_ex
    .imme(imme_num),
    .rdata_a(rdata_a),
    .rdata_b(rdata_b),
    .greater_than(greater_than),
    .equal_branch(equal_branch),
    .bgtz_sig(bgtz_sig),
    .zero_sig(zero_sig),
    .jc_instaddress(jc_instaddress)
);

opcode_control opcode_control(
    .opcode(opcode),
    .RegDst(RegDst),
    .Branch(Branch),
    .MemRead(MemRead),
    .MemtoReg(MemtoReg),
    .ALUOp(ALUOp),
    .MemWrite(MemWrite),
    .ALUSrc(ALUSrc),
    .RegWrite(RegWrite),
    .Jump(Jump),
    .equal_branch(equal_branch),
    .store_pc(store_pc),
    .lui_sig(lui_sig),
    .greater_than(greater_than)
);

regs regs(
    .clk(clk),
    .rst(rst),
    .rreg_a(rreg_a),
    .rreg_b(rreg_b),
    .wreg(mem_wreg),
    .wdata(mem_wdata),
    .RegWrite(mem_RegWrite),
    .rdata_a(rdata_a),
    .rdata_b(rdata_b),
    .inst_address(ex_cur_instaddress),
    .store_pc(ex_store_pc)
);

pre_alu pre_alu(
    .ex_rdata_a(ex_rdata_a),
    .ex_rdata_b(ex_rdata_b),
    .mem_wb_dout(mem_wdata),
    .control_rdata_a(control_rdata_a),
    .control_rdata_b(control_rdata_b),
    .rdata_a(alu_rdata_a),
    .rdata_b(alu_rdata_b)
);

alu alu(
    .data_a(alu_rdata_a),
    .data_b(alu_rdata_b),
    .imme(ex_imme_num),
    .ALUSrc(ex_ALUSrc),
    .alu_control(alu_control_sig),
    //.zero_sig(ALU_zerotag),
    .alu_result(alu_result),
    .unsigned_num(unsigned_num),
    .equal_branch(ex_equal_branch),
    .shamt(ex_shamt)
    //.greater_than(ex_greater_than),
    //.bgtz_sig(bgtz_sig)
);

alu_control alu_control(
    .func(ex_func),
    .ALUOp(ex_ALUOp),
    .opcode(ex_opcode),
    .alu_control(alu_control_sig)
);

pre_mem pre_mem(
    .opcode(mem_opcode),
    .mem_sel(mem_sel)
);

mem mem(
    .clk(clk),
    .alu_result(mem_alu_result),
    .din(mem_rdata_b),            //���ԼĴ����ѵĵڶ�����������
    .MemWrite(mem_MemWrite),
    .MemRead(mem_MemRead),
    .MemtoReg(mem_MemtoReg),
    .dout(mem_wdata),
    .mem_sel(mem_sel),
    .lui_sig(mem_lui_sig),
    //.mem_wreg(mem_wreg),
    //.mem_RegWrite(mem_RegWrite),
    //.wb_RegWrite(wb_RegWrite),
    //.wb_wreg(wb_wreg),
    .imme(mem_imme_num)            //����id�׶ε�������
);

redirect redirect(
    .ex_Rs(ex_Rs),
    .ex_Rt(ex_Rt),
    .mem_wb_wreg(mem_wreg),
    .mem_wb_RegWrite(mem_RegWrite),
    .control_rdata_a(control_rdata_a),
    .control_rdata_b(control_rdata_b)
);

endmodule