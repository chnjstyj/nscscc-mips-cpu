module inst_rom(                 //ָ��Ĵ���
    input clk,
    input rom_clk,
    input [31:0] inst_address,
    input ce,
    output reg read_ce,
    output [31:0] irom_addr,
    input [31:0] rom_inst,
    input rfin_c,
    input rfin_d,
    /*
    input [15:0] rdata_a,
    input [15:0] rdata_b,
    output [31:0] rom_addr,
    output rom_ce,
    output we,
    output oe,
    output reg [31:0] inst 
    */
);

//reg [31:0] inst_rom[0:1023];      //4kb��reg
//reg read_ce;
//reg [31:0] address;
assign irom_addr = {inst_address[31:2],2'b00};

//wire [15:0] data_a;
//wire [15:0] data_b;
//wire rfin;

//initial $readmemh( "F:\inst_rom.data", inst_rom );

/*
always @(*) begin
    if(ce == 1'b0) begin 
        inst <= 32'h00000000;
    end 
    else begin 
        inst <= inst_rom[inst_address[11:2]];
    end 
end */

//���ڴ�
always @(*) begin 
    if(ce == 1'b0) begin
        inst <= 32'h00000000;
        read_ce <= 1'b0;
    end 
    else begin 
        read_ce <= 1'b1;
        if(rfin_c && rfin_d) inst <= rom_inst;
        else inst <= inst;
    end
end
/*
mips ���ֽ�Ѱַ������ָ���ַҪ/2�������λ��ȡ��
��log2(1024) = 10,����ֻȡǰ10λ��
*/
/*
irom_read irom_read_a(
    .clk(rom_clk),
    .rst(rst),
    .read_ce(read_ce),
    .address(address),
    .dout(rdata_a),
    .data(data_a),
    .rfin(rfin),
    .ce(rom_ce),
    .we(we),
    .oe(oe)
);

irom_read irom_read_b(
    .clk(rom_clk),
    .rst(rst),
    .read_ce(read_ce),
    .address(address),
    .dout(rdata_b),
    .data(data_b),
    .rfin(rfin),
    .ce(rom_ce),
    .we(we),
    .oe(oe)
);
*/

endmodule  